module test_coordinator(); endmodule