module task (
    input  [15:0] a,        // 第一个16位操作数
    input  [15:0] b,        // 第二个16位操作数  
    input         cin,      // 输入进位
    output [15:0] sum,      // 16位和
    output        cout      // 输出进位
);

// 定义内部信号
wire [15:0] g;  // 进位生成信号
wire [15:0] p;  // 进位传播信号
wire [15:0] carry;  // 中间进位信号

// 计算每个位的进位生成 (G) 和进位传播 (P)
genvar i;
generate
    for (i = 0; i < 16; i = i + 1) begin : gen_g_p
        assign g[i] = a[i] & b[i];
        assign p[i] = a[i] ^ b[i];
    end
endgenerate

// 初始化第一个进位
assign carry[0] = cin;

// 递归计算进位
generate
    for (i = 1; i < 16; i = i + 1) begin : gen_carry
        assign carry[i] = g[i-1] | (p[i-1] & carry[i-1]);
    end
endgenerate

// 计算和
generate
    for (i = 0; i < 16; i = i + 1) begin : gen_sum
        assign sum[i] = p[i] ^ carry[i];
    end
endgenerate

// 最终进位输出
assign cout = carry[15];

endmodule