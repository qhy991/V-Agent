module simple_8bit_adder (
    input  [7:0] a,         // 第一个8位操作数
    input  [7:0] b,         // 第二个8位操作数
    input        cin,       // 输入进位
    output wire [7:0] sum,  // 8位和
    output wire       cout  // 输出进位
);

    // 内部信号声明
    wire [7:0] carry;

    // 第一位加法器（最低位）
    full_adder fa0 (
        .a(a[0]),
        .b(b[0]),
        .cin(cin),
        .sum(sum[0]),
        .cout(carry[0])
    );

    // 其余7位加法器
    generate
        for (integer i = 1; i < 8; i = i + 1) begin : adder_loop
            full_adder fa (
                .a(a[i]),
                .b(b[i]),
                .cin(carry[i-1]),
                .sum(sum[i]),
                .cout(carry[i])
            );
        end
    endgenerate

    // 输出进位是最高位的进位
    assign cout = carry[7];

endmodule

// 全加器子模块
module full_adder (
    input  a,
    input  b,
    input  cin,
    output sum,
    output cout
);

    // 计算和
    assign sum = a ^ b ^ cin;

    // 计算进位
    assign cout = (a & b) | (a & cin) | (b & cin);

endmodule