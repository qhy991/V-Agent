module test_tool_call(); endmodule