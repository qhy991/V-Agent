// 临时依赖文件
module temp_module; endmodule