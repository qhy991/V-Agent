// Quick test file
module quick_test();
endmodule