module test_path(); endmodule