// Test file for function calling
module test();
endmodule