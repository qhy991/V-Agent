module alu;
endmodule;