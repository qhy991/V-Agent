module simple_8bit_adder (
// Full adder module definition
module full_adder (
endmodule
endmodule