// Performance test file 0
module test_0();
endmodule