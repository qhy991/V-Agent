module counter_8bit;
  // Module description: 8-bit counter with synchronous reset, enable control, and overflow flag
endmodule;