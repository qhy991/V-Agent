module simple_8bit_adder (
endmodule