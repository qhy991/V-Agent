module test2(); endmodule