module empty_module();
endmodule