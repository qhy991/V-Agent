module task (
endmodule