// Performance test file 1
module test_1();
endmodule