module simple_8bit_adder (
module full_adder (
endmodule
endmodule