module counter_with_comments (
    input      clk,     // 时钟信号，上升沿触发
    input      reset,   // 同步复位信号，高电平有效
    input      enable,  // 计数使能信号，高电平允许计数
    output reg [7:0] count  // 当前8位计数值输出
);

// ============================================================================
// 模块功能描述：
// 该模块实现一个8位同步复位、使能控制的递增计数器。
// 在时钟上升沿，当enable信号为高电平时，计数器递增；
// 当reset信号为高电平时，计数器同步清零。
// ============================================================================
// 端口说明：
// - clk: 主时钟信号，上升沿触发计数操作
// - reset: 同步复位信号，高电平有效，优先于enable
// - enable: 使能信号，控制是否允许计数递增
// - count: 8位输出寄存器，表示当前计数值
// ============================================================================

// 内部逻辑实现
always @(posedge clk) begin : counter_proc
    // 在时钟上升沿执行操作
    if (reset) begin
        // 复位条件成立时，将计数器清零
        count <= 8'h00;
    end else if (enable) begin
        // 使能信号有效时，计数器递增
        count <= count + 1;
    end
    // 如果reset为低且enable为低，保持当前计数值不变
end

endmodule