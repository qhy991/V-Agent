module test_enhanced(); endmodule