
module test();
    initial begin
        $display("Hello from test module!");
        $finish;
    end
endmodule
