module alu_32bit (
endmodule