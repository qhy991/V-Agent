// Performance test file 2
module test_2();
endmodule