module test(); endmodule