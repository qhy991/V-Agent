module adder_4bit (
endmodule