module unknown_module();
endmodule