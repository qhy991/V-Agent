module carry_lookahead_adder_16bit (
endmodule